%RC circuit

R1 1 0 1
R2 2 0 1
R3 3 0 1
R4 1 2 1
R5 2 3 1

I1 1 0 1

.op
.end
